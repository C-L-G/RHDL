module  XXXX  //head comment
/*
    body comment
*/
/*
parameter PPP

endparameter

interface III

endinterface

localparam LLL

endlocalparamr
*/
endmodule:
