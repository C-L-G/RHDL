module  XXXX

endmodule
