module  XXXX

interface IIII
endinterface

endmodule
